module main

import tinyid

fn main() {
	println(tinyid.new(12))
}
